-- EASE/HDL begin --------------------------------------------------------------
-- 
-- Architecture 'behavior' of entity 'div_freq'.
-- 
--------------------------------------------------------------------------------
-- 
-- Copy of the interface declaration:
-- 
--   port (
--     clk     : in     std_logic;
--     div     : in     std_logic_vector(15 downto 0);
--     freq    : out    std_logic;
--     reset_n : in     std_logic);
-- 
-- EASE/HDL end ----------------------------------------------------------------

architecture behavior of div_freq is

begin

end architecture behavior ; -- of div_freq

