-- EASE/HDL begin --------------------------------------------------------------
-- 
-- Architecture 'behavior' of entity 'counter_sec'.
-- 
--------------------------------------------------------------------------------
-- 
-- Copy of the interface declaration:
-- 
--   port (
--     clk     : in     std_logic;
--     freq    : in     std_logic;
--     reset_n : in     std_logic;
--     s_pulse : out    std_logic);
-- 
-- EASE/HDL end ----------------------------------------------------------------

architecture behavior of counter_sec is

begin

end architecture behavior ; -- of counter_sec

