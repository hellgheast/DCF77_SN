-- EASE/HDL begin --------------------------------------------------------------
-- 
-- Architecture 'behavioral' of entity 'counter_ms_oveflow'.
-- 
--------------------------------------------------------------------------------
-- 
-- Copy of the interface declaration:
-- 
--   port (
--     clk                : in     std_logic;
--     freq               : in     std_logic;
--     reset_n            : in     std_logic;
--     rising_edge_dcf_77 : in     std_logic;
--     sec_overflow       : out    std_logic);
-- 
-- EASE/HDL end ----------------------------------------------------------------

architecture behavioral of counter_ms_oveflow is

begin

end architecture behavioral ; -- of counter_ms_oveflow

