-- EASE/HDL begin --------------------------------------------------------------
-- 
-- Architecture 'behavioral' of entity 'rising_edge_dectection'.
-- 
--------------------------------------------------------------------------------
-- 
-- Copy of the interface declaration:
-- 
-- EASE/HDL end ----------------------------------------------------------------

architecture behavioral of rising_edge_dectection is

begin

end architecture behavioral ; -- of rising_edge_dectection

