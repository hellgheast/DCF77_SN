-- EASE/HDL begin --------------------------------------------------------------
-- 
-- Architecture 'behavior' of entity 'DecodeStateMachine'.
-- 
--------------------------------------------------------------------------------
-- 
-- Copy of the interface declaration:
-- 
-- EASE/HDL end ----------------------------------------------------------------

architecture behavior of DecodeStateMachine is

begin

end architecture behavior ; -- of DecodeStateMachine

