-- EASE/HDL begin --------------------------------------------------------------
-- 
-- Architecture 'behavior' of entity 'frame_register'.
-- 
--------------------------------------------------------------------------------
-- 
-- Copy of the interface declaration:
-- 
--   port (
--     RBG         : in     std_logic_vector(2 downto 0);
--     bit         : in     std_logic;
--     bit_count   : in     std_logic_vector(5 downto 0);
--     clk         : in     std_logic;
--     reg_dmonth  : out    std_logic_vector(6 downto 0);
--     reg_dweek   : out    std_logic_vector(2 downto 0);
--     reg_flags   : out    std_logic_vector(3 downto 0);
--     reg_hours   : out    std_logic_vector(5 downto 0);
--     reg_minutes : out    std_logic_vector(6 downto 0);
--     reg_month   : out    std_logic_vector(5 downto 0);
--     reg_status  : out    std_logic_vector(7 downto 0);
--     reg_year    : out    std_logic_vector(7 downto 0);
--     reset_n     : in     std_logic;
--     start       : in     std_logic;
--     stop        : in     std_logic);
-- 
-- EASE/HDL end ----------------------------------------------------------------

architecture behavior of frame_register is

begin

end architecture behavior ; -- of frame_register

