-- EASE/HDL begin --------------------------------------------------------------
-- 
-- Architecture 'behavior' of entity 'reg_mem_dcf77'.
-- 
--------------------------------------------------------------------------------
-- 
-- Copy of the interface declaration:
-- 
--   port (
--     Adress      : in     std_logic_vector(3 downto 0);
--     chip_select : in     std_logic;
--     clk         : in     std_logic;
--     data_in     : in     std_logic_vector(7 downto 0);
--     data_out    : out    std_logic_vector(7 downto 0);
--     prescaler   : out    std_logic_vector(15 downto 0);
--     read        : in     std_logic;
--     reg_dmonth  : in     std_logic_vector(6 downto 0);
--     reg_dweek   : in     std_logic_vector(2 downto 0);
--     reg_flags   : in     std_logic_vector(3 downto 0);
--     reg_hours   : in     std_logic_vector(5 downto 0);
--     reg_minutes : in     std_logic_vector(6 downto 0);
--     reg_month   : in     std_logic_vector(5 downto 0);
--     reg_status  : in     std_logic_vector(7 downto 0);
--     reg_year    : in     std_logic_vector(7 downto 0);
--     reset_n     : in     std_logic;
--     write       : in     std_logic);
-- 
-- EASE/HDL end ----------------------------------------------------------------

architecture behavior of reg_mem_dcf77 is

begin

end architecture behavior ; -- of reg_mem_dcf77

