-- EASE/HDL begin --------------------------------------------------------------
-- 
-- Architecture 'behavior' of entity 'decode_RBG'.
-- 
--------------------------------------------------------------------------------
-- 
-- Copy of the interface declaration:
-- 
--   port (
--     RBG       : out    std_logic_vector(2 downto 0);
--     bit_count : in     std_logic_vector(5 downto 0);
--     start     : in     std_logic;
--     stop      : in     std_logic);
-- 
-- EASE/HDL end ----------------------------------------------------------------

architecture behavior of decode_RBG is

begin     

if bit_count 

end architecture behavior ; -- of decode_RBG

